tt06Endo REACTION { initialState = tt06Endo; }
tt06Endo SINGLECELL {
  method = BetterTT06;
  Vm = -85.851589919619585 mV;
  Ca_SR = 3.3928054282480442 uM;
  Ca_i = 0.00010226128163141762 uM;
  Ca_ss = 0.00018549989458331147 uM;
  K_i = 137.60835983603508 mM;
  Na_i = 9.6613086409123454 mM;
  R_prime = 0.98937816635116493 1;
  Xr1 = -1.0801626442798633e-05 1;
  Xr2 = 0.47878870593482692 1;
  Xs = 0.0031059009148968696 1;
  d = 1.0039861458801012e-05 1;
  f = 0.97765812635714333 1;
  f2 = 0.99958790918010709 1;
  fCass = 0.99997517999320673 1;
  h = 0.75954312065793239 1;
  j = 0.75924727373539103 1;
  m = 0.0013261154521225097 1;
  r = 5.271986789650334e-06 1;
  s = 0.64641686415579114 1;
}
