tt06Mid REACTION { initialState = tt06Mid; }
tt06Mid SINGLECELL {
  method = BetterTT06;
  Vm = -85.70769745705914 mV;
  Ca_SR = 4.1316479299519395 uM;
  Ca_i = 0.00011550656128389796 uM;
  Ca_ss = 0.00020820387700369328 uM;
  K_i = 137.64493896206264 mM;
  Na_i = 9.4957688259918296 mM;
  R_prime = 0.98765885854718849 1;
  Xr1 = -8.3202368746061153e-07 1;
  Xr2 = 0.47728915796059557 1;
  Xs = 0.0032245967822579244 1;
  d = 1.0308124465673115e-05 1;
  f = 0.96043927822410402 1;
  f2 = 0.99936384991278049 1;
  fCass = 0.99996431717350387 1;
  h = 0.7558015594316615 1;
  j = 0.75515365697618897 1;
  m = 0.0013756261848726907 1;
  r = 5.2764699914834664e-06 1;
  s = 0.99995080955034976 1;
}
